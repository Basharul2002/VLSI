module my_not(input wire A,
              output wire Y)
  not(Y,A)
endmodule
