module or(input wire A, B
           output wire Y)
  or(Y, A,B)
endmodule
        
