module xor(input wire A, B,
           output wire Y);
  xor(Y, A, B);
endmodule
