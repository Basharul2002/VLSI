module nor(input wire A, B,
            output wire Y);
  nor(Y, A,B);
endmodule
