module nand(input wire A, B,
            output wire Y);
  nand(Y, A,B);
endmodule
