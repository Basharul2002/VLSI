module and(input wire A, B
           output wire Y)
  and(Y, A,B)
endmodule
        
