module xnor(input wire A, B,
            output wire Y);
  xnor(Y, A,B);
endmodule
